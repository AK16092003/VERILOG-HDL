`timescale 1ns / 1ns
`include "division.v"

module division_tb;
	
reg [2:0] D;
reg [1:0] V;

wire [2:0] Q;
wire [1:0] R;
wire Z;

division uut(D,V,Q,R,Z);
initial
	$monitor($time,"ns  D = %b ,V = %b ,Q = %b ,R = %b ,Z = %b " , D,V,Q,R,Z);
initial begin
	$dumpfile("division_tb.vcd");
	$dumpvars(0,division_tb);
	
	D[2] = 0;D[1] = 0;D[0] = 0;
	V[1] = 0;V[0] = 0;
	#2;
	D[2] = 0;D[1] = 0;D[0] = 0;
	V[1] = 0;V[0] = 1;
	#2;
	D[2] = 0;D[1] = 0;D[0] = 0;
	V[1] = 1;V[0] = 0;
	#2;
	D[2] = 0;D[1] = 0;D[0] = 0;
	V[1] = 1;V[0] = 1;
	#2;
	D[2] = 0;D[1] = 0;D[0] = 1;
	V[1] = 0;V[0] = 0;
	#2;
	D[2] = 0;D[1] = 0;D[0] = 1;
	V[1] = 0;V[0] = 1;
	#2;
	D[2] = 0;D[1] = 0;D[0] = 1;
	V[1] = 1;V[0] = 0;
	#2;
	D[2] = 0;D[1] = 0;D[0] = 1;
	V[1] = 1;V[0] = 1;
	#2;
	D[2] = 0;D[1] = 1;D[0] = 0;
	V[1] = 0;V[0] = 0;
	#2;
	D[2] = 0;D[1] = 1;D[0] = 0;
	V[1] = 0;V[0] = 1;
	#2;
	D[2] = 0;D[1] = 1;D[0] = 0;
	V[1] = 1;V[0] = 0;
	#2;
	D[2] = 0;D[1] = 1;D[0] = 0;
	V[1] = 1;V[0] = 1;
	#2;
	D[2] = 0;D[1] = 1;D[0] = 1;
	V[1] = 0;V[0] = 0;
	#2;
	D[2] = 0;D[1] = 1;D[0] = 1;
	V[1] = 0;V[0] = 1;
	#2;
	D[2] = 0;D[1] = 1;D[0] = 1;
	V[1] = 1;V[0] = 0;
	#2;
	D[2] = 0;D[1] = 1;D[0] = 1;
	V[1] = 1;V[0] = 1;
	#2;
	D[2] = 1;D[1] = 0;D[0] = 0;
	V[1] = 0;V[0] = 0;
	#2;
	D[2] = 1;D[1] = 0;D[0] = 0;
	V[1] = 0;V[0] = 1;
	#2;
	D[2] = 1;D[1] = 0;D[0] = 0;
	V[1] = 1;V[0] = 0;
	#2;
	D[2] = 1;D[1] = 0;D[0] = 0;
	V[1] = 1;V[0] = 1;
	#2;
	D[2] = 1;D[1] = 0;D[0] = 1;
	V[1] = 0;V[0] = 0;
	#2;
	D[2] = 1;D[1] = 0;D[0] = 1;
	V[1] = 0;V[0] = 1;
	#2;
	D[2] = 1;D[1] = 0;D[0] = 1;
	V[1] = 1;V[0] = 0;
	#2;
	D[2] = 1;D[1] = 0;D[0] = 1;
	V[1] = 1;V[0] = 1;
	#2;
	D[2] = 1;D[1] = 1;D[0] = 0;
	V[1] = 0;V[0] = 0;
	#2;
	D[2] = 1;D[1] = 1;D[0] = 0;
	V[1] = 0;V[0] = 1;
	#2;
	D[2] = 1;D[1] = 1;D[0] = 0;
	V[1] = 1;V[0] = 0;
	#2;
	D[2] = 1;D[1] = 1;D[0] = 0;
	V[1] = 1;V[0] = 1;
	#2;
	D[2] = 1;D[1] = 1;D[0] = 1;
	V[1] = 0;V[0] = 0;
	#2;
	D[2] = 1;D[1] = 1;D[0] = 1;
	V[1] = 0;V[0] = 1;
	#2;
	D[2] = 1;D[1] = 1;D[0] = 1;
	V[1] = 1;V[0] = 0;
	#2;
	D[2] = 1;D[1] = 1;D[0] = 1;
	V[1] = 1;V[0] = 1;
	#2;
	$display("Test completed ");	
end
endmodule